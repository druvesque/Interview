// Q. Design a sequence detector for 101011 (overlapping)?
//
// Q. Write an assertion in SystemVerilog such that if a then 
//    b should be high for the next 2 clock cycles.
//
// Q. Describe different types of arrays in SystemVerilog.
//
// Q. What is your approach to ensure quality in a product? 
//
// Q. Explain always block in verilog and always_comb, always_ff
//    & always_latch in SystemVerilog with the help of code.
