// Q1. 
