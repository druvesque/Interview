// Q. I2C Project Explanation
//
//    - In my project, I implemented a complete I2C communication system 
//      in Verilog by designing both the master and slave controllers.
//      I created FSM to check start and stop conditions, handle address
//      transmission, data transfer and acknowledge cycles. 
//
//    - I also implemented clock generation logic for SCL and open-drain
//      Style SDA control. On the slave side, I designed the address decoding
//      And data response logic. 
