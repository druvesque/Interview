// Q. Explain FIFO and what different types of FIFOs are there?
//
//    - FIFO is a buffer that stores data such that the first data written
//      is the first data read.
//
//    - Synchronous FIFO
//      Same clock for read and write.
