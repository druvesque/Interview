// Q1. Is UVM independent of SystemVerilog
//
//     - No, UVM is built on SystemVerilog and hence you cannot
//       run UVM with any tool that does not support SystemVerilog.
